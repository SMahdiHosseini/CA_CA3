module DP(input[2:0] AluOperation,input[1:0] PCSrc,input[1:0] AluSrcB,input rst,clk,PcSrc,link,RegDst,RegWrite,AluSrcA,
	IRWrite,MemWrite,MemRead,MemtoReg,PCWrite,PCWriteCond,branch,output[5:0] func,output[5:0] opcode);
		
	
endmodule
